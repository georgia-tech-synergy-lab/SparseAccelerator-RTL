../../accelerator/data_control/output_control.sv