../../accelerator/vegeta_top.sv