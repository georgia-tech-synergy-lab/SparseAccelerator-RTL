../../accelerator/data_control/vegeta_control.sv