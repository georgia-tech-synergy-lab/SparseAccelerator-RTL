../../accelerator/compute/vegeta_pu.sv