../../accelerator/compute/vegeta_compute_top.sv