../../accelerator/arithmetic/fp32_adder.sv