../../accelerator/arithmetic/bf16_mult.sv