../../accelerator/data_control/accumulation_control.sv