../../accelerator/data_control/activation_control.sv