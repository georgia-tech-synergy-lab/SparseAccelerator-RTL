../../accelerator/compute/vegeta_mac.sv