../../accelerator/arithmetic/general_adder.sv