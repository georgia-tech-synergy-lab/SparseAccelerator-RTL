../../accelerator/compute/vegeta_pe.sv