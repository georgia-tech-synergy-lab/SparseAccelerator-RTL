../../accelerator/testbenches/vegeta_top_tb/vegeta_top_tb.sv