../../accelerator/compute/adder_tree.sv