../../accelerator/data_control/weight_control.sv