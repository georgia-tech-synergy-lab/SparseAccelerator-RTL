../../accelerator/arithmetic/general_multiplier.sv