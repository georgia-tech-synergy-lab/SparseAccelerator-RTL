../../accelerator/memory/L1_buffer.sv