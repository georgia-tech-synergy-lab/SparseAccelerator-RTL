../../accelerator/memory/L1_buffer_independent_write.sv